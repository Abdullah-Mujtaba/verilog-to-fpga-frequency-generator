`timescale 1ns / 1ps
`define S6_TO_U8(x) {x, 2'b00}

module DDS(
    input clk,
    input reset,
    input [9:0] ftw,    
    output reg [7:0] sin_wave
);

reg [9:0] rotation;
reg [9:0] index;

always @(posedge clk) begin
    if (reset) begin
        rotation <= 0;
        index <= 0;
    end
    else begin
        rotation <= rotation + ftw; 
        index <= rotation;
    end
end

always @(*) begin
    case (index)
        10'h000: sin_wave = `S6_TO_U8(6'h1F);
        10'h001: sin_wave = `S6_TO_U8(6'h1F);
        10'h002: sin_wave = `S6_TO_U8(6'h1F);
        10'h003: sin_wave = `S6_TO_U8(6'h20);
        10'h004: sin_wave = `S6_TO_U8(6'h20);
        10'h005: sin_wave = `S6_TO_U8(6'h20);
        10'h006: sin_wave = `S6_TO_U8(6'h20);
        10'h007: sin_wave = `S6_TO_U8(6'h20);
        10'h008: sin_wave = `S6_TO_U8(6'h21);
        10'h009: sin_wave = `S6_TO_U8(6'h21);
        10'h00A: sin_wave = `S6_TO_U8(6'h21);
        10'h00B: sin_wave = `S6_TO_U8(6'h21);
        10'h00C: sin_wave = `S6_TO_U8(6'h21);
        10'h00D: sin_wave = `S6_TO_U8(6'h22);
        10'h00E: sin_wave = `S6_TO_U8(6'h22);
        10'h00F: sin_wave = `S6_TO_U8(6'h22);
        10'h010: sin_wave = `S6_TO_U8(6'h22);
        10'h011: sin_wave = `S6_TO_U8(6'h22);
        10'h012: sin_wave = `S6_TO_U8(6'h22);
        10'h013: sin_wave = `S6_TO_U8(6'h23);
        10'h014: sin_wave = `S6_TO_U8(6'h23);
        10'h015: sin_wave = `S6_TO_U8(6'h23);
        10'h016: sin_wave = `S6_TO_U8(6'h23);
        10'h017: sin_wave = `S6_TO_U8(6'h23);
        10'h018: sin_wave = `S6_TO_U8(6'h24);
        10'h019: sin_wave = `S6_TO_U8(6'h24);
        10'h01A: sin_wave = `S6_TO_U8(6'h24);
        10'h01B: sin_wave = `S6_TO_U8(6'h24);
        10'h01C: sin_wave = `S6_TO_U8(6'h24);
        10'h01D: sin_wave = `S6_TO_U8(6'h25);
        10'h01E: sin_wave = `S6_TO_U8(6'h25);
        10'h01F: sin_wave = `S6_TO_U8(6'h25);
        10'h020: sin_wave = `S6_TO_U8(6'h25);
        10'h021: sin_wave = `S6_TO_U8(6'h25);
        10'h022: sin_wave = `S6_TO_U8(6'h26);
        10'h023: sin_wave = `S6_TO_U8(6'h26);
        10'h024: sin_wave = `S6_TO_U8(6'h26);
        10'h025: sin_wave = `S6_TO_U8(6'h26);
        10'h026: sin_wave = `S6_TO_U8(6'h26);
        10'h027: sin_wave = `S6_TO_U8(6'h26);
        10'h028: sin_wave = `S6_TO_U8(6'h27);
        10'h029: sin_wave = `S6_TO_U8(6'h27);
        10'h02A: sin_wave = `S6_TO_U8(6'h27);
        10'h02B: sin_wave = `S6_TO_U8(6'h27);
        10'h02C: sin_wave = `S6_TO_U8(6'h27);
        10'h02D: sin_wave = `S6_TO_U8(6'h28);
        10'h02E: sin_wave = `S6_TO_U8(6'h28);
        10'h02F: sin_wave = `S6_TO_U8(6'h28);
        10'h030: sin_wave = `S6_TO_U8(6'h28);
        10'h031: sin_wave = `S6_TO_U8(6'h28);
        10'h032: sin_wave = `S6_TO_U8(6'h29);
        10'h033: sin_wave = `S6_TO_U8(6'h29);
        10'h034: sin_wave = `S6_TO_U8(6'h29);
        10'h035: sin_wave = `S6_TO_U8(6'h29);
        10'h036: sin_wave = `S6_TO_U8(6'h29);
        10'h037: sin_wave = `S6_TO_U8(6'h29);
        10'h038: sin_wave = `S6_TO_U8(6'h2A);
        10'h039: sin_wave = `S6_TO_U8(6'h2A);
        10'h03A: sin_wave = `S6_TO_U8(6'h2A);
        10'h03B: sin_wave = `S6_TO_U8(6'h2A);
        10'h03C: sin_wave = `S6_TO_U8(6'h2A);
        10'h03D: sin_wave = `S6_TO_U8(6'h2B);
        10'h03E: sin_wave = `S6_TO_U8(6'h2B);
        10'h03F: sin_wave = `S6_TO_U8(6'h2B);
        10'h040: sin_wave = `S6_TO_U8(6'h2B);
        10'h041: sin_wave = `S6_TO_U8(6'h2B);
        10'h042: sin_wave = `S6_TO_U8(6'h2B);
        10'h043: sin_wave = `S6_TO_U8(6'h2C);
        10'h044: sin_wave = `S6_TO_U8(6'h2C);
        10'h045: sin_wave = `S6_TO_U8(6'h2C);
        10'h046: sin_wave = `S6_TO_U8(6'h2C);
        10'h047: sin_wave = `S6_TO_U8(6'h2C);
        10'h048: sin_wave = `S6_TO_U8(6'h2C);
        10'h049: sin_wave = `S6_TO_U8(6'h2D);
        10'h04A: sin_wave = `S6_TO_U8(6'h2D);
        10'h04B: sin_wave = `S6_TO_U8(6'h2D);
        10'h04C: sin_wave = `S6_TO_U8(6'h2D);
        10'h04D: sin_wave = `S6_TO_U8(6'h2D);
        10'h04E: sin_wave = `S6_TO_U8(6'h2E);
        10'h04F: sin_wave = `S6_TO_U8(6'h2E);
        10'h050: sin_wave = `S6_TO_U8(6'h2E);
        10'h051: sin_wave = `S6_TO_U8(6'h2E);
        10'h052: sin_wave = `S6_TO_U8(6'h2E);
        10'h053: sin_wave = `S6_TO_U8(6'h2E);
        10'h054: sin_wave = `S6_TO_U8(6'h2F);
        10'h055: sin_wave = `S6_TO_U8(6'h2F);
        10'h056: sin_wave = `S6_TO_U8(6'h2F);
        10'h057: sin_wave = `S6_TO_U8(6'h2F);
        10'h058: sin_wave = `S6_TO_U8(6'h2F);
        10'h059: sin_wave = `S6_TO_U8(6'h2F);
        10'h05A: sin_wave = `S6_TO_U8(6'h30);
        10'h05B: sin_wave = `S6_TO_U8(6'h30);
        10'h05C: sin_wave = `S6_TO_U8(6'h30);
        10'h05D: sin_wave = `S6_TO_U8(6'h30);
        10'h05E: sin_wave = `S6_TO_U8(6'h30);
        10'h05F: sin_wave = `S6_TO_U8(6'h30);
        10'h060: sin_wave = `S6_TO_U8(6'h31);
        10'h061: sin_wave = `S6_TO_U8(6'h31);
        10'h062: sin_wave = `S6_TO_U8(6'h31);
        10'h063: sin_wave = `S6_TO_U8(6'h31);
        10'h064: sin_wave = `S6_TO_U8(6'h31);
        10'h065: sin_wave = `S6_TO_U8(6'h31);
        10'h066: sin_wave = `S6_TO_U8(6'h31);
        10'h067: sin_wave = `S6_TO_U8(6'h32);
        10'h068: sin_wave = `S6_TO_U8(6'h32);
        10'h069: sin_wave = `S6_TO_U8(6'h32);
        10'h06A: sin_wave = `S6_TO_U8(6'h32);
        10'h06B: sin_wave = `S6_TO_U8(6'h32);
        10'h06C: sin_wave = `S6_TO_U8(6'h32);
        10'h06D: sin_wave = `S6_TO_U8(6'h33);
        10'h06E: sin_wave = `S6_TO_U8(6'h33);
        10'h06F: sin_wave = `S6_TO_U8(6'h33);
        10'h070: sin_wave = `S6_TO_U8(6'h33);
        10'h071: sin_wave = `S6_TO_U8(6'h33);
        10'h072: sin_wave = `S6_TO_U8(6'h33);
        10'h073: sin_wave = `S6_TO_U8(6'h33);
        10'h074: sin_wave = `S6_TO_U8(6'h34);
        10'h075: sin_wave = `S6_TO_U8(6'h34);
        10'h076: sin_wave = `S6_TO_U8(6'h34);
        10'h077: sin_wave = `S6_TO_U8(6'h34);
        10'h078: sin_wave = `S6_TO_U8(6'h34);
        10'h079: sin_wave = `S6_TO_U8(6'h34);
        10'h07A: sin_wave = `S6_TO_U8(6'h34);
        10'h07B: sin_wave = `S6_TO_U8(6'h35);
        10'h07C: sin_wave = `S6_TO_U8(6'h35);
        10'h07D: sin_wave = `S6_TO_U8(6'h35);
        10'h07E: sin_wave = `S6_TO_U8(6'h35);
        10'h07F: sin_wave = `S6_TO_U8(6'h35);
        10'h080: sin_wave = `S6_TO_U8(6'h35);
        10'h081: sin_wave = `S6_TO_U8(6'h35);
        10'h082: sin_wave = `S6_TO_U8(6'h36);
        10'h083: sin_wave = `S6_TO_U8(6'h36);
        10'h084: sin_wave = `S6_TO_U8(6'h36);
        10'h085: sin_wave = `S6_TO_U8(6'h36);
        10'h086: sin_wave = `S6_TO_U8(6'h36);
        10'h087: sin_wave = `S6_TO_U8(6'h36);
        10'h088: sin_wave = `S6_TO_U8(6'h36);
        10'h089: sin_wave = `S6_TO_U8(6'h36);
        10'h08A: sin_wave = `S6_TO_U8(6'h37);
        10'h08B: sin_wave = `S6_TO_U8(6'h37);
        10'h08C: sin_wave = `S6_TO_U8(6'h37);
        10'h08D: sin_wave = `S6_TO_U8(6'h37);
        10'h08E: sin_wave = `S6_TO_U8(6'h37);
        10'h08F: sin_wave = `S6_TO_U8(6'h37);
        10'h090: sin_wave = `S6_TO_U8(6'h37);
        10'h091: sin_wave = `S6_TO_U8(6'h37);
        10'h092: sin_wave = `S6_TO_U8(6'h38);
        10'h093: sin_wave = `S6_TO_U8(6'h38);
        10'h094: sin_wave = `S6_TO_U8(6'h38);
        10'h095: sin_wave = `S6_TO_U8(6'h38);
        10'h096: sin_wave = `S6_TO_U8(6'h38);
        10'h097: sin_wave = `S6_TO_U8(6'h38);
        10'h098: sin_wave = `S6_TO_U8(6'h38);
        10'h099: sin_wave = `S6_TO_U8(6'h38);
        10'h09A: sin_wave = `S6_TO_U8(6'h39);
        10'h09B: sin_wave = `S6_TO_U8(6'h39);
        10'h09C: sin_wave = `S6_TO_U8(6'h39);
        10'h09D: sin_wave = `S6_TO_U8(6'h39);
        10'h09E: sin_wave = `S6_TO_U8(6'h39);
        10'h09F: sin_wave = `S6_TO_U8(6'h39);
        10'h0A0: sin_wave = `S6_TO_U8(6'h39);
        10'h0A1: sin_wave = `S6_TO_U8(6'h39);
        10'h0A2: sin_wave = `S6_TO_U8(6'h39);
        10'h0A3: sin_wave = `S6_TO_U8(6'h3A);
        10'h0A4: sin_wave = `S6_TO_U8(6'h3A);
        10'h0A5: sin_wave = `S6_TO_U8(6'h3A);
        10'h0A6: sin_wave = `S6_TO_U8(6'h3A);
        10'h0A7: sin_wave = `S6_TO_U8(6'h3A);
        10'h0A8: sin_wave = `S6_TO_U8(6'h3A);
        10'h0A9: sin_wave = `S6_TO_U8(6'h3A);
        10'h0AA: sin_wave = `S6_TO_U8(6'h3A);
        10'h0AB: sin_wave = `S6_TO_U8(6'h3A);
        10'h0AC: sin_wave = `S6_TO_U8(6'h3A);
        10'h0AD: sin_wave = `S6_TO_U8(6'h3B);
        10'h0AE: sin_wave = `S6_TO_U8(6'h3B);
        10'h0AF: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B0: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B1: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B2: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B3: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B4: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B5: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B6: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B7: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B8: sin_wave = `S6_TO_U8(6'h3B);
        10'h0B9: sin_wave = `S6_TO_U8(6'h3C);
        10'h0BA: sin_wave = `S6_TO_U8(6'h3C);
        10'h0BB: sin_wave = `S6_TO_U8(6'h3C);
        10'h0BC: sin_wave = `S6_TO_U8(6'h3C);
        10'h0BD: sin_wave = `S6_TO_U8(6'h3C);
        10'h0BE: sin_wave = `S6_TO_U8(6'h3C);
        10'h0BF: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C0: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C1: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C2: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C3: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C4: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C5: sin_wave = `S6_TO_U8(6'h3C);
        10'h0C6: sin_wave = `S6_TO_U8(6'h3D);
        10'h0C7: sin_wave = `S6_TO_U8(6'h3D);
        10'h0C8: sin_wave = `S6_TO_U8(6'h3D);
        10'h0C9: sin_wave = `S6_TO_U8(6'h3D);
        10'h0CA: sin_wave = `S6_TO_U8(6'h3D);
        10'h0CB: sin_wave = `S6_TO_U8(6'h3D);
        10'h0CC: sin_wave = `S6_TO_U8(6'h3D);
        10'h0CD: sin_wave = `S6_TO_U8(6'h3D);
        10'h0CE: sin_wave = `S6_TO_U8(6'h3D);
        10'h0CF: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D0: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D1: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D2: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D3: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D4: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D5: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D6: sin_wave = `S6_TO_U8(6'h3D);
        10'h0D7: sin_wave = `S6_TO_U8(6'h3E);
        10'h0D8: sin_wave = `S6_TO_U8(6'h3E);
        10'h0D9: sin_wave = `S6_TO_U8(6'h3E);
        10'h0DA: sin_wave = `S6_TO_U8(6'h3E);
        10'h0DB: sin_wave = `S6_TO_U8(6'h3E);
        10'h0DC: sin_wave = `S6_TO_U8(6'h3E);
        10'h0DD: sin_wave = `S6_TO_U8(6'h3E);
        10'h0DE: sin_wave = `S6_TO_U8(6'h3E);
        10'h0DF: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E0: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E1: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E2: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E3: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E4: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E5: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E6: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E7: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E8: sin_wave = `S6_TO_U8(6'h3E);
        10'h0E9: sin_wave = `S6_TO_U8(6'h3E);
        10'h0EA: sin_wave = `S6_TO_U8(6'h3E);
        10'h0EB: sin_wave = `S6_TO_U8(6'h3E);
        10'h0EC: sin_wave = `S6_TO_U8(6'h3E);
        10'h0ED: sin_wave = `S6_TO_U8(6'h3E);
        10'h0EE: sin_wave = `S6_TO_U8(6'h3E);
        10'h0EF: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F0: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F1: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F2: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F3: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F4: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F5: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F6: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F7: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F8: sin_wave = `S6_TO_U8(6'h3E);
        10'h0F9: sin_wave = `S6_TO_U8(6'h3E);
        10'h0FA: sin_wave = `S6_TO_U8(6'h3E);
        10'h0FB: sin_wave = `S6_TO_U8(6'h3E);
        10'h0FC: sin_wave = `S6_TO_U8(6'h3E);
        10'h0FD: sin_wave = `S6_TO_U8(6'h3E);
        10'h0FE: sin_wave = `S6_TO_U8(6'h3E);
        10'h0FF: sin_wave = `S6_TO_U8(6'h3E);
        10'h100: sin_wave = `S6_TO_U8(6'h3F);
        10'h101: sin_wave = `S6_TO_U8(6'h3E);
        10'h102: sin_wave = `S6_TO_U8(6'h3E);
        10'h103: sin_wave = `S6_TO_U8(6'h3E);
        10'h104: sin_wave = `S6_TO_U8(6'h3E);
        10'h105: sin_wave = `S6_TO_U8(6'h3E);
        10'h106: sin_wave = `S6_TO_U8(6'h3E);
        10'h107: sin_wave = `S6_TO_U8(6'h3E);
        10'h108: sin_wave = `S6_TO_U8(6'h3E);
        10'h109: sin_wave = `S6_TO_U8(6'h3E);
        10'h10A: sin_wave = `S6_TO_U8(6'h3E);
        10'h10B: sin_wave = `S6_TO_U8(6'h3E);
        10'h10C: sin_wave = `S6_TO_U8(6'h3E);
        10'h10D: sin_wave = `S6_TO_U8(6'h3E);
        10'h10E: sin_wave = `S6_TO_U8(6'h3E);
        10'h10F: sin_wave = `S6_TO_U8(6'h3E);
        10'h110: sin_wave = `S6_TO_U8(6'h3E);
        10'h111: sin_wave = `S6_TO_U8(6'h3E);
        10'h112: sin_wave = `S6_TO_U8(6'h3E);
        10'h113: sin_wave = `S6_TO_U8(6'h3E);
        10'h114: sin_wave = `S6_TO_U8(6'h3E);
        10'h115: sin_wave = `S6_TO_U8(6'h3E);
        10'h116: sin_wave = `S6_TO_U8(6'h3E);
        10'h117: sin_wave = `S6_TO_U8(6'h3E);
        10'h118: sin_wave = `S6_TO_U8(6'h3E);
        10'h119: sin_wave = `S6_TO_U8(6'h3E);
        10'h11A: sin_wave = `S6_TO_U8(6'h3E);
        10'h11B: sin_wave = `S6_TO_U8(6'h3E);
        10'h11C: sin_wave = `S6_TO_U8(6'h3E);
        10'h11D: sin_wave = `S6_TO_U8(6'h3E);
        10'h11E: sin_wave = `S6_TO_U8(6'h3E);
        10'h11F: sin_wave = `S6_TO_U8(6'h3E);
        10'h120: sin_wave = `S6_TO_U8(6'h3E);
        10'h121: sin_wave = `S6_TO_U8(6'h3E);
        10'h122: sin_wave = `S6_TO_U8(6'h3E);
        10'h123: sin_wave = `S6_TO_U8(6'h3E);
        10'h124: sin_wave = `S6_TO_U8(6'h3E);
        10'h125: sin_wave = `S6_TO_U8(6'h3E);
        10'h126: sin_wave = `S6_TO_U8(6'h3E);
        10'h127: sin_wave = `S6_TO_U8(6'h3E);
        10'h128: sin_wave = `S6_TO_U8(6'h3E);
        10'h129: sin_wave = `S6_TO_U8(6'h3E);
        10'h12A: sin_wave = `S6_TO_U8(6'h3D);
        10'h12B: sin_wave = `S6_TO_U8(6'h3D);
        10'h12C: sin_wave = `S6_TO_U8(6'h3D);
        10'h12D: sin_wave = `S6_TO_U8(6'h3D);
        10'h12E: sin_wave = `S6_TO_U8(6'h3D);
        10'h12F: sin_wave = `S6_TO_U8(6'h3D);
        10'h130: sin_wave = `S6_TO_U8(6'h3D);
        10'h131: sin_wave = `S6_TO_U8(6'h3D);
        10'h132: sin_wave = `S6_TO_U8(6'h3D);
        10'h133: sin_wave = `S6_TO_U8(6'h3D);
        10'h134: sin_wave = `S6_TO_U8(6'h3D);
        10'h135: sin_wave = `S6_TO_U8(6'h3D);
        10'h136: sin_wave = `S6_TO_U8(6'h3D);
        10'h137: sin_wave = `S6_TO_U8(6'h3D);
        10'h138: sin_wave = `S6_TO_U8(6'h3D);
        10'h139: sin_wave = `S6_TO_U8(6'h3D);
        10'h13A: sin_wave = `S6_TO_U8(6'h3D);
        10'h13B: sin_wave = `S6_TO_U8(6'h3C);
        10'h13C: sin_wave = `S6_TO_U8(6'h3C);
        10'h13D: sin_wave = `S6_TO_U8(6'h3C);
        10'h13E: sin_wave = `S6_TO_U8(6'h3C);
        10'h13F: sin_wave = `S6_TO_U8(6'h3C);
        10'h140: sin_wave = `S6_TO_U8(6'h3C);
        10'h141: sin_wave = `S6_TO_U8(6'h3C);
        10'h142: sin_wave = `S6_TO_U8(6'h3C);
        10'h143: sin_wave = `S6_TO_U8(6'h3C);
        10'h144: sin_wave = `S6_TO_U8(6'h3C);
        10'h145: sin_wave = `S6_TO_U8(6'h3C);
        10'h146: sin_wave = `S6_TO_U8(6'h3C);
        10'h147: sin_wave = `S6_TO_U8(6'h3C);
        10'h148: sin_wave = `S6_TO_U8(6'h3B);
        10'h149: sin_wave = `S6_TO_U8(6'h3B);
        10'h14A: sin_wave = `S6_TO_U8(6'h3B);
        10'h14B: sin_wave = `S6_TO_U8(6'h3B);
        10'h14C: sin_wave = `S6_TO_U8(6'h3B);
        10'h14D: sin_wave = `S6_TO_U8(6'h3B);
        10'h14E: sin_wave = `S6_TO_U8(6'h3B);
        10'h14F: sin_wave = `S6_TO_U8(6'h3B);
        10'h150: sin_wave = `S6_TO_U8(6'h3B);
        10'h151: sin_wave = `S6_TO_U8(6'h3B);
        10'h152: sin_wave = `S6_TO_U8(6'h3B);
        10'h153: sin_wave = `S6_TO_U8(6'h3B);
        10'h154: sin_wave = `S6_TO_U8(6'h3A);
        10'h155: sin_wave = `S6_TO_U8(6'h3A);
        10'h156: sin_wave = `S6_TO_U8(6'h3A);
        10'h157: sin_wave = `S6_TO_U8(6'h3A);
        10'h158: sin_wave = `S6_TO_U8(6'h3A);
        10'h159: sin_wave = `S6_TO_U8(6'h3A);
        10'h15A: sin_wave = `S6_TO_U8(6'h3A);
        10'h15B: sin_wave = `S6_TO_U8(6'h3A);
        10'h15C: sin_wave = `S6_TO_U8(6'h3A);
        10'h15D: sin_wave = `S6_TO_U8(6'h3A);
        10'h15E: sin_wave = `S6_TO_U8(6'h39);
        10'h15F: sin_wave = `S6_TO_U8(6'h39);
        10'h160: sin_wave = `S6_TO_U8(6'h39);
        10'h161: sin_wave = `S6_TO_U8(6'h39);
        10'h162: sin_wave = `S6_TO_U8(6'h39);
        10'h163: sin_wave = `S6_TO_U8(6'h39);
        10'h164: sin_wave = `S6_TO_U8(6'h39);
        10'h165: sin_wave = `S6_TO_U8(6'h39);
        10'h166: sin_wave = `S6_TO_U8(6'h39);
        10'h167: sin_wave = `S6_TO_U8(6'h38);
        10'h168: sin_wave = `S6_TO_U8(6'h38);
        10'h169: sin_wave = `S6_TO_U8(6'h38);
        10'h16A: sin_wave = `S6_TO_U8(6'h38);
        10'h16B: sin_wave = `S6_TO_U8(6'h38);
        10'h16C: sin_wave = `S6_TO_U8(6'h38);
        10'h16D: sin_wave = `S6_TO_U8(6'h38);
        10'h16E: sin_wave = `S6_TO_U8(6'h38);
        10'h16F: sin_wave = `S6_TO_U8(6'h37);
        10'h170: sin_wave = `S6_TO_U8(6'h37);
        10'h171: sin_wave = `S6_TO_U8(6'h37);
        10'h172: sin_wave = `S6_TO_U8(6'h37);
        10'h173: sin_wave = `S6_TO_U8(6'h37);
        10'h174: sin_wave = `S6_TO_U8(6'h37);
        10'h175: sin_wave = `S6_TO_U8(6'h37);
        10'h176: sin_wave = `S6_TO_U8(6'h37);
        10'h177: sin_wave = `S6_TO_U8(6'h36);
        10'h178: sin_wave = `S6_TO_U8(6'h36);
        10'h179: sin_wave = `S6_TO_U8(6'h36);
        10'h17A: sin_wave = `S6_TO_U8(6'h36);
        10'h17B: sin_wave = `S6_TO_U8(6'h36);
        10'h17C: sin_wave = `S6_TO_U8(6'h36);
        10'h17D: sin_wave = `S6_TO_U8(6'h36);
        10'h17E: sin_wave = `S6_TO_U8(6'h36);
        10'h17F: sin_wave = `S6_TO_U8(6'h35);
        10'h180: sin_wave = `S6_TO_U8(6'h35);
        10'h181: sin_wave = `S6_TO_U8(6'h35);
        10'h182: sin_wave = `S6_TO_U8(6'h35);
        10'h183: sin_wave = `S6_TO_U8(6'h35);
        10'h184: sin_wave = `S6_TO_U8(6'h35);
        10'h185: sin_wave = `S6_TO_U8(6'h35);
        10'h186: sin_wave = `S6_TO_U8(6'h34);
        10'h187: sin_wave = `S6_TO_U8(6'h34);
        10'h188: sin_wave = `S6_TO_U8(6'h34);
        10'h189: sin_wave = `S6_TO_U8(6'h34);
        10'h18A: sin_wave = `S6_TO_U8(6'h34);
        10'h18B: sin_wave = `S6_TO_U8(6'h34);
        10'h18C: sin_wave = `S6_TO_U8(6'h34);
        10'h18D: sin_wave = `S6_TO_U8(6'h33);
        10'h18E: sin_wave = `S6_TO_U8(6'h33);
        10'h18F: sin_wave = `S6_TO_U8(6'h33);
        10'h190: sin_wave = `S6_TO_U8(6'h33);
        10'h191: sin_wave = `S6_TO_U8(6'h33);
        10'h192: sin_wave = `S6_TO_U8(6'h33);
        10'h193: sin_wave = `S6_TO_U8(6'h33);
        10'h194: sin_wave = `S6_TO_U8(6'h32);
        10'h195: sin_wave = `S6_TO_U8(6'h32);
        10'h196: sin_wave = `S6_TO_U8(6'h32);
        10'h197: sin_wave = `S6_TO_U8(6'h32);
        10'h198: sin_wave = `S6_TO_U8(6'h32);
        10'h199: sin_wave = `S6_TO_U8(6'h32);
        10'h19A: sin_wave = `S6_TO_U8(6'h31);
        10'h19B: sin_wave = `S6_TO_U8(6'h31);
        10'h19C: sin_wave = `S6_TO_U8(6'h31);
        10'h19D: sin_wave = `S6_TO_U8(6'h31);
        10'h19E: sin_wave = `S6_TO_U8(6'h31);
        10'h19F: sin_wave = `S6_TO_U8(6'h31);
        10'h1A0: sin_wave = `S6_TO_U8(6'h31);
        10'h1A1: sin_wave = `S6_TO_U8(6'h30);
        10'h1A2: sin_wave = `S6_TO_U8(6'h30);
        10'h1A3: sin_wave = `S6_TO_U8(6'h30);
        10'h1A4: sin_wave = `S6_TO_U8(6'h30);
        10'h1A5: sin_wave = `S6_TO_U8(6'h30);
        10'h1A6: sin_wave = `S6_TO_U8(6'h30);
        10'h1A7: sin_wave = `S6_TO_U8(6'h2F);
        10'h1A8: sin_wave = `S6_TO_U8(6'h2F);
        10'h1A9: sin_wave = `S6_TO_U8(6'h2F);
        10'h1AA: sin_wave = `S6_TO_U8(6'h2F);
        10'h1AB: sin_wave = `S6_TO_U8(6'h2F);
        10'h1AC: sin_wave = `S6_TO_U8(6'h2F);
        10'h1AD: sin_wave = `S6_TO_U8(6'h2E);
        10'h1AE: sin_wave = `S6_TO_U8(6'h2E);
        10'h1AF: sin_wave = `S6_TO_U8(6'h2E);
        10'h1B0: sin_wave = `S6_TO_U8(6'h2E);
        10'h1B1: sin_wave = `S6_TO_U8(6'h2E);
        10'h1B2: sin_wave = `S6_TO_U8(6'h2E);
        10'h1B3: sin_wave = `S6_TO_U8(6'h2D);
        10'h1B4: sin_wave = `S6_TO_U8(6'h2D);
        10'h1B5: sin_wave = `S6_TO_U8(6'h2D);
        10'h1B6: sin_wave = `S6_TO_U8(6'h2D);
        10'h1B7: sin_wave = `S6_TO_U8(6'h2D);
        10'h1B8: sin_wave = `S6_TO_U8(6'h2C);
        10'h1B9: sin_wave = `S6_TO_U8(6'h2C);
        10'h1BA: sin_wave = `S6_TO_U8(6'h2C);
        10'h1BB: sin_wave = `S6_TO_U8(6'h2C);
        10'h1BC: sin_wave = `S6_TO_U8(6'h2C);
        10'h1BD: sin_wave = `S6_TO_U8(6'h2C);
        10'h1BE: sin_wave = `S6_TO_U8(6'h2B);
        10'h1BF: sin_wave = `S6_TO_U8(6'h2B);
        10'h1C0: sin_wave = `S6_TO_U8(6'h2B);
        10'h1C1: sin_wave = `S6_TO_U8(6'h2B);
        10'h1C2: sin_wave = `S6_TO_U8(6'h2B);
        10'h1C3: sin_wave = `S6_TO_U8(6'h2B);
        10'h1C4: sin_wave = `S6_TO_U8(6'h2A);
        10'h1C5: sin_wave = `S6_TO_U8(6'h2A);
        10'h1C6: sin_wave = `S6_TO_U8(6'h2A);
        10'h1C7: sin_wave = `S6_TO_U8(6'h2A);
        10'h1C8: sin_wave = `S6_TO_U8(6'h2A);
        10'h1C9: sin_wave = `S6_TO_U8(6'h29);
        10'h1CA: sin_wave = `S6_TO_U8(6'h29);
        10'h1CB: sin_wave = `S6_TO_U8(6'h29);
        10'h1CC: sin_wave = `S6_TO_U8(6'h29);
        10'h1CD: sin_wave = `S6_TO_U8(6'h29);
        10'h1CE: sin_wave = `S6_TO_U8(6'h29);
        10'h1CF: sin_wave = `S6_TO_U8(6'h28);
        10'h1D0: sin_wave = `S6_TO_U8(6'h28);
        10'h1D1: sin_wave = `S6_TO_U8(6'h28);
        10'h1D2: sin_wave = `S6_TO_U8(6'h28);
        10'h1D3: sin_wave = `S6_TO_U8(6'h28);
        10'h1D4: sin_wave = `S6_TO_U8(6'h27);
        10'h1D5: sin_wave = `S6_TO_U8(6'h27);
        10'h1D6: sin_wave = `S6_TO_U8(6'h27);
        10'h1D7: sin_wave = `S6_TO_U8(6'h27);
        10'h1D8: sin_wave = `S6_TO_U8(6'h27);
        10'h1D9: sin_wave = `S6_TO_U8(6'h26);
        10'h1DA: sin_wave = `S6_TO_U8(6'h26);
        10'h1DB: sin_wave = `S6_TO_U8(6'h26);
        10'h1DC: sin_wave = `S6_TO_U8(6'h26);
        10'h1DD: sin_wave = `S6_TO_U8(6'h26);
        10'h1DE: sin_wave = `S6_TO_U8(6'h26);
        10'h1DF: sin_wave = `S6_TO_U8(6'h25);
        10'h1E0: sin_wave = `S6_TO_U8(6'h25);
        10'h1E1: sin_wave = `S6_TO_U8(6'h25);
        10'h1E2: sin_wave = `S6_TO_U8(6'h25);
        10'h1E3: sin_wave = `S6_TO_U8(6'h25);
        10'h1E4: sin_wave = `S6_TO_U8(6'h24);
        10'h1E5: sin_wave = `S6_TO_U8(6'h24);
        10'h1E6: sin_wave = `S6_TO_U8(6'h24);
        10'h1E7: sin_wave = `S6_TO_U8(6'h24);
        10'h1E8: sin_wave = `S6_TO_U8(6'h24);
        10'h1E9: sin_wave = `S6_TO_U8(6'h23);
        10'h1EA: sin_wave = `S6_TO_U8(6'h23);
        10'h1EB: sin_wave = `S6_TO_U8(6'h23);
        10'h1EC: sin_wave = `S6_TO_U8(6'h23);
        10'h1ED: sin_wave = `S6_TO_U8(6'h23);
        10'h1EE: sin_wave = `S6_TO_U8(6'h22);
        10'h1EF: sin_wave = `S6_TO_U8(6'h22);
        10'h1F0: sin_wave = `S6_TO_U8(6'h22);
        10'h1F1: sin_wave = `S6_TO_U8(6'h22);
        10'h1F2: sin_wave = `S6_TO_U8(6'h22);
        10'h1F3: sin_wave = `S6_TO_U8(6'h22);
        10'h1F4: sin_wave = `S6_TO_U8(6'h21);
        10'h1F5: sin_wave = `S6_TO_U8(6'h21);
        10'h1F6: sin_wave = `S6_TO_U8(6'h21);
        10'h1F7: sin_wave = `S6_TO_U8(6'h21);
        10'h1F8: sin_wave = `S6_TO_U8(6'h21);
        10'h1F9: sin_wave = `S6_TO_U8(6'h20);
        10'h1FA: sin_wave = `S6_TO_U8(6'h20);
        10'h1FB: sin_wave = `S6_TO_U8(6'h20);
        10'h1FC: sin_wave = `S6_TO_U8(6'h20);
        10'h1FD: sin_wave = `S6_TO_U8(6'h20);
        10'h1FE: sin_wave = `S6_TO_U8(6'h1F);
        10'h1FF: sin_wave = `S6_TO_U8(6'h1F);
        10'h200: sin_wave = `S6_TO_U8(6'h1F);
        10'h201: sin_wave = `S6_TO_U8(6'h1F);
        10'h202: sin_wave = `S6_TO_U8(6'h1F);
        10'h203: sin_wave = `S6_TO_U8(6'h1E);
        10'h204: sin_wave = `S6_TO_U8(6'h1E);
        10'h205: sin_wave = `S6_TO_U8(6'h1E);
        10'h206: sin_wave = `S6_TO_U8(6'h1E);
        10'h207: sin_wave = `S6_TO_U8(6'h1E);
        10'h208: sin_wave = `S6_TO_U8(6'h1D);
        10'h209: sin_wave = `S6_TO_U8(6'h1D);
        10'h20A: sin_wave = `S6_TO_U8(6'h1D);
        10'h20B: sin_wave = `S6_TO_U8(6'h1D);
        10'h20C: sin_wave = `S6_TO_U8(6'h1D);
        10'h20D: sin_wave = `S6_TO_U8(6'h1C);
        10'h20E: sin_wave = `S6_TO_U8(6'h1C);
        10'h20F: sin_wave = `S6_TO_U8(6'h1C);
        10'h210: sin_wave = `S6_TO_U8(6'h1C);
        10'h211: sin_wave = `S6_TO_U8(6'h1C);
        10'h212: sin_wave = `S6_TO_U8(6'h1C);
        10'h213: sin_wave = `S6_TO_U8(6'h1B);
        10'h214: sin_wave = `S6_TO_U8(6'h1B);
        10'h215: sin_wave = `S6_TO_U8(6'h1B);
        10'h216: sin_wave = `S6_TO_U8(6'h1B);
        10'h217: sin_wave = `S6_TO_U8(6'h1B);
        10'h218: sin_wave = `S6_TO_U8(6'h1A);
        10'h219: sin_wave = `S6_TO_U8(6'h1A);
        10'h21A: sin_wave = `S6_TO_U8(6'h1A);
        10'h21B: sin_wave = `S6_TO_U8(6'h1A);
        10'h21C: sin_wave = `S6_TO_U8(6'h1A);
        10'h21D: sin_wave = `S6_TO_U8(6'h19);
        10'h21E: sin_wave = `S6_TO_U8(6'h19);
        10'h21F: sin_wave = `S6_TO_U8(6'h19);
        10'h220: sin_wave = `S6_TO_U8(6'h19);
        10'h221: sin_wave = `S6_TO_U8(6'h19);
        10'h222: sin_wave = `S6_TO_U8(6'h18);
        10'h223: sin_wave = `S6_TO_U8(6'h18);
        10'h224: sin_wave = `S6_TO_U8(6'h18);
        10'h225: sin_wave = `S6_TO_U8(6'h18);
        10'h226: sin_wave = `S6_TO_U8(6'h18);
        10'h227: sin_wave = `S6_TO_U8(6'h18);
        10'h228: sin_wave = `S6_TO_U8(6'h17);
        10'h229: sin_wave = `S6_TO_U8(6'h17);
        10'h22A: sin_wave = `S6_TO_U8(6'h17);
        10'h22B: sin_wave = `S6_TO_U8(6'h17);
        10'h22C: sin_wave = `S6_TO_U8(6'h17);
        10'h22D: sin_wave = `S6_TO_U8(6'h16);
        10'h22E: sin_wave = `S6_TO_U8(6'h16);
        10'h22F: sin_wave = `S6_TO_U8(6'h16);
        10'h230: sin_wave = `S6_TO_U8(6'h16);
        10'h231: sin_wave = `S6_TO_U8(6'h16);
        10'h232: sin_wave = `S6_TO_U8(6'h15);
        10'h233: sin_wave = `S6_TO_U8(6'h15);
        10'h234: sin_wave = `S6_TO_U8(6'h15);
        10'h235: sin_wave = `S6_TO_U8(6'h15);
        10'h236: sin_wave = `S6_TO_U8(6'h15);
        10'h237: sin_wave = `S6_TO_U8(6'h15);
        10'h238: sin_wave = `S6_TO_U8(6'h14);
        10'h239: sin_wave = `S6_TO_U8(6'h14);
        10'h23A: sin_wave = `S6_TO_U8(6'h14);
        10'h23B: sin_wave = `S6_TO_U8(6'h14);
        10'h23C: sin_wave = `S6_TO_U8(6'h14);
        10'h23D: sin_wave = `S6_TO_U8(6'h13);
        10'h23E: sin_wave = `S6_TO_U8(6'h13);
        10'h23F: sin_wave = `S6_TO_U8(6'h13);
        10'h240: sin_wave = `S6_TO_U8(6'h13);
        10'h241: sin_wave = `S6_TO_U8(6'h13);
        10'h242: sin_wave = `S6_TO_U8(6'h13);
        10'h243: sin_wave = `S6_TO_U8(6'h12);
        10'h244: sin_wave = `S6_TO_U8(6'h12);
        10'h245: sin_wave = `S6_TO_U8(6'h12);
        10'h246: sin_wave = `S6_TO_U8(6'h12);
        10'h247: sin_wave = `S6_TO_U8(6'h12);
        10'h248: sin_wave = `S6_TO_U8(6'h12);
        10'h249: sin_wave = `S6_TO_U8(6'h11);
        10'h24A: sin_wave = `S6_TO_U8(6'h11);
        10'h24B: sin_wave = `S6_TO_U8(6'h11);
        10'h24C: sin_wave = `S6_TO_U8(6'h11);
        10'h24D: sin_wave = `S6_TO_U8(6'h11);
        10'h24E: sin_wave = `S6_TO_U8(6'h10);
        10'h24F: sin_wave = `S6_TO_U8(6'h10);
        10'h250: sin_wave = `S6_TO_U8(6'h10);
        10'h251: sin_wave = `S6_TO_U8(6'h10);
        10'h252: sin_wave = `S6_TO_U8(6'h10);
        10'h253: sin_wave = `S6_TO_U8(6'h10);
        10'h254: sin_wave = `S6_TO_U8(6'h0F);
        10'h255: sin_wave = `S6_TO_U8(6'h0F);
        10'h256: sin_wave = `S6_TO_U8(6'h0F);
        10'h257: sin_wave = `S6_TO_U8(6'h0F);
        10'h258: sin_wave = `S6_TO_U8(6'h0F);
        10'h259: sin_wave = `S6_TO_U8(6'h0F);
        10'h25A: sin_wave = `S6_TO_U8(6'h0E);
        10'h25B: sin_wave = `S6_TO_U8(6'h0E);
        10'h25C: sin_wave = `S6_TO_U8(6'h0E);
        10'h25D: sin_wave = `S6_TO_U8(6'h0E);
        10'h25E: sin_wave = `S6_TO_U8(6'h0E);
        10'h25F: sin_wave = `S6_TO_U8(6'h0E);
        10'h260: sin_wave = `S6_TO_U8(6'h0D);
        10'h261: sin_wave = `S6_TO_U8(6'h0D);
        10'h262: sin_wave = `S6_TO_U8(6'h0D);
        10'h263: sin_wave = `S6_TO_U8(6'h0D);
        10'h264: sin_wave = `S6_TO_U8(6'h0D);
        10'h265: sin_wave = `S6_TO_U8(6'h0D);
        10'h266: sin_wave = `S6_TO_U8(6'h0D);
        10'h267: sin_wave = `S6_TO_U8(6'h0C);
        10'h268: sin_wave = `S6_TO_U8(6'h0C);
        10'h269: sin_wave = `S6_TO_U8(6'h0C);
        10'h26A: sin_wave = `S6_TO_U8(6'h0C);
        10'h26B: sin_wave = `S6_TO_U8(6'h0C);
        10'h26C: sin_wave = `S6_TO_U8(6'h0C);
        10'h26D: sin_wave = `S6_TO_U8(6'h0B);
        10'h26E: sin_wave = `S6_TO_U8(6'h0B);
        10'h26F: sin_wave = `S6_TO_U8(6'h0B);
        10'h270: sin_wave = `S6_TO_U8(6'h0B);
        10'h271: sin_wave = `S6_TO_U8(6'h0B);
        10'h272: sin_wave = `S6_TO_U8(6'h0B);
        10'h273: sin_wave = `S6_TO_U8(6'h0B);
        10'h274: sin_wave = `S6_TO_U8(6'h0A);
        10'h275: sin_wave = `S6_TO_U8(6'h0A);
        10'h276: sin_wave = `S6_TO_U8(6'h0A);
        10'h277: sin_wave = `S6_TO_U8(6'h0A);
        10'h278: sin_wave = `S6_TO_U8(6'h0A);
        10'h279: sin_wave = `S6_TO_U8(6'h0A);
        10'h27A: sin_wave = `S6_TO_U8(6'h0A);
        10'h27B: sin_wave = `S6_TO_U8(6'h09);
        10'h27C: sin_wave = `S6_TO_U8(6'h09);
        10'h27D: sin_wave = `S6_TO_U8(6'h09);
        10'h27E: sin_wave = `S6_TO_U8(6'h09);
        10'h27F: sin_wave = `S6_TO_U8(6'h09);
        10'h280: sin_wave = `S6_TO_U8(6'h09);
        10'h281: sin_wave = `S6_TO_U8(6'h09);
        10'h282: sin_wave = `S6_TO_U8(6'h08);
        10'h283: sin_wave = `S6_TO_U8(6'h08);
        10'h284: sin_wave = `S6_TO_U8(6'h08);
        10'h285: sin_wave = `S6_TO_U8(6'h08);
        10'h286: sin_wave = `S6_TO_U8(6'h08);
        10'h287: sin_wave = `S6_TO_U8(6'h08);
        10'h288: sin_wave = `S6_TO_U8(6'h08);
        10'h289: sin_wave = `S6_TO_U8(6'h08);
        10'h28A: sin_wave = `S6_TO_U8(6'h07);
        10'h28B: sin_wave = `S6_TO_U8(6'h07);
        10'h28C: sin_wave = `S6_TO_U8(6'h07);
        10'h28D: sin_wave = `S6_TO_U8(6'h07);
        10'h28E: sin_wave = `S6_TO_U8(6'h07);
        10'h28F: sin_wave = `S6_TO_U8(6'h07);
        10'h290: sin_wave = `S6_TO_U8(6'h07);
        10'h291: sin_wave = `S6_TO_U8(6'h07);
        10'h292: sin_wave = `S6_TO_U8(6'h06);
        10'h293: sin_wave = `S6_TO_U8(6'h06);
        10'h294: sin_wave = `S6_TO_U8(6'h06);
        10'h295: sin_wave = `S6_TO_U8(6'h06);
        10'h296: sin_wave = `S6_TO_U8(6'h06);
        10'h297: sin_wave = `S6_TO_U8(6'h06);
        10'h298: sin_wave = `S6_TO_U8(6'h06);
        10'h299: sin_wave = `S6_TO_U8(6'h06);
        10'h29A: sin_wave = `S6_TO_U8(6'h05);
        10'h29B: sin_wave = `S6_TO_U8(6'h05);
        10'h29C: sin_wave = `S6_TO_U8(6'h05);
        10'h29D: sin_wave = `S6_TO_U8(6'h05);
        10'h29E: sin_wave = `S6_TO_U8(6'h05);
        10'h29F: sin_wave = `S6_TO_U8(6'h05);
        10'h2A0: sin_wave = `S6_TO_U8(6'h05);
        10'h2A1: sin_wave = `S6_TO_U8(6'h05);
        10'h2A2: sin_wave = `S6_TO_U8(6'h05);
        10'h2A3: sin_wave = `S6_TO_U8(6'h04);
        10'h2A4: sin_wave = `S6_TO_U8(6'h04);
        10'h2A5: sin_wave = `S6_TO_U8(6'h04);
        10'h2A6: sin_wave = `S6_TO_U8(6'h04);
        10'h2A7: sin_wave = `S6_TO_U8(6'h04);
        10'h2A8: sin_wave = `S6_TO_U8(6'h04);
        10'h2A9: sin_wave = `S6_TO_U8(6'h04);
        10'h2AA: sin_wave = `S6_TO_U8(6'h04);
        10'h2AB: sin_wave = `S6_TO_U8(6'h04);
        10'h2AC: sin_wave = `S6_TO_U8(6'h04);
        10'h2AD: sin_wave = `S6_TO_U8(6'h03);
        10'h2AE: sin_wave = `S6_TO_U8(6'h03);
        10'h2AF: sin_wave = `S6_TO_U8(6'h03);
        10'h2B0: sin_wave = `S6_TO_U8(6'h03);
        10'h2B1: sin_wave = `S6_TO_U8(6'h03);
        10'h2B2: sin_wave = `S6_TO_U8(6'h03);
        10'h2B3: sin_wave = `S6_TO_U8(6'h03);
        10'h2B4: sin_wave = `S6_TO_U8(6'h03);
        10'h2B5: sin_wave = `S6_TO_U8(6'h03);
        10'h2B6: sin_wave = `S6_TO_U8(6'h03);
        10'h2B7: sin_wave = `S6_TO_U8(6'h03);
        10'h2B8: sin_wave = `S6_TO_U8(6'h03);
        10'h2B9: sin_wave = `S6_TO_U8(6'h02);
        10'h2BA: sin_wave = `S6_TO_U8(6'h02);
        10'h2BB: sin_wave = `S6_TO_U8(6'h02);
        10'h2BC: sin_wave = `S6_TO_U8(6'h02);
        10'h2BD: sin_wave = `S6_TO_U8(6'h02);
        10'h2BE: sin_wave = `S6_TO_U8(6'h02);
        10'h2BF: sin_wave = `S6_TO_U8(6'h02);
        10'h2C0: sin_wave = `S6_TO_U8(6'h02);
        10'h2C1: sin_wave = `S6_TO_U8(6'h02);
        10'h2C2: sin_wave = `S6_TO_U8(6'h02);
        10'h2C3: sin_wave = `S6_TO_U8(6'h02);
        10'h2C4: sin_wave = `S6_TO_U8(6'h02);
        10'h2C5: sin_wave = `S6_TO_U8(6'h02);
        10'h2C6: sin_wave = `S6_TO_U8(6'h01);
        10'h2C7: sin_wave = `S6_TO_U8(6'h01);
        10'h2C8: sin_wave = `S6_TO_U8(6'h01);
        10'h2C9: sin_wave = `S6_TO_U8(6'h01);
        10'h2CA: sin_wave = `S6_TO_U8(6'h01);
        10'h2CB: sin_wave = `S6_TO_U8(6'h01);
        10'h2CC: sin_wave = `S6_TO_U8(6'h01);
        10'h2CD: sin_wave = `S6_TO_U8(6'h01);
        10'h2CE: sin_wave = `S6_TO_U8(6'h01);
        10'h2CF: sin_wave = `S6_TO_U8(6'h01);
        10'h2D0: sin_wave = `S6_TO_U8(6'h01);
        10'h2D1: sin_wave = `S6_TO_U8(6'h01);
        10'h2D2: sin_wave = `S6_TO_U8(6'h01);
        10'h2D3: sin_wave = `S6_TO_U8(6'h01);
        10'h2D4: sin_wave = `S6_TO_U8(6'h01);
        10'h2D5: sin_wave = `S6_TO_U8(6'h01);
        10'h2D6: sin_wave = `S6_TO_U8(6'h01);
        10'h2D7: sin_wave = `S6_TO_U8(6'h00);
        10'h2D8: sin_wave = `S6_TO_U8(6'h00);
        10'h2D9: sin_wave = `S6_TO_U8(6'h00);
        10'h2DA: sin_wave = `S6_TO_U8(6'h00);
        10'h2DB: sin_wave = `S6_TO_U8(6'h00);
        10'h2DC: sin_wave = `S6_TO_U8(6'h00);
        10'h2DD: sin_wave = `S6_TO_U8(6'h00);
        10'h2DE: sin_wave = `S6_TO_U8(6'h00);
        10'h2DF: sin_wave = `S6_TO_U8(6'h00);
        10'h2E0: sin_wave = `S6_TO_U8(6'h00);
        10'h2E1: sin_wave = `S6_TO_U8(6'h00);
        10'h2E2: sin_wave = `S6_TO_U8(6'h00);
        10'h2E3: sin_wave = `S6_TO_U8(6'h00);
        10'h2E4: sin_wave = `S6_TO_U8(6'h00);
        10'h2E5: sin_wave = `S6_TO_U8(6'h00);
        10'h2E6: sin_wave = `S6_TO_U8(6'h00);
        10'h2E7: sin_wave = `S6_TO_U8(6'h00);
        10'h2E8: sin_wave = `S6_TO_U8(6'h00);
        10'h2E9: sin_wave = `S6_TO_U8(6'h00);
        10'h2EA: sin_wave = `S6_TO_U8(6'h00);
        10'h2EB: sin_wave = `S6_TO_U8(6'h00);
        10'h2EC: sin_wave = `S6_TO_U8(6'h00);
        10'h2ED: sin_wave = `S6_TO_U8(6'h00);
        10'h2EE: sin_wave = `S6_TO_U8(6'h00);
        10'h2EF: sin_wave = `S6_TO_U8(6'h00);
        10'h2F0: sin_wave = `S6_TO_U8(6'h00);
        10'h2F1: sin_wave = `S6_TO_U8(6'h00);
        10'h2F2: sin_wave = `S6_TO_U8(6'h00);
        10'h2F3: sin_wave = `S6_TO_U8(6'h00);
        10'h2F4: sin_wave = `S6_TO_U8(6'h00);
        10'h2F5: sin_wave = `S6_TO_U8(6'h00);
        10'h2F6: sin_wave = `S6_TO_U8(6'h00);
        10'h2F7: sin_wave = `S6_TO_U8(6'h00);
        10'h2F8: sin_wave = `S6_TO_U8(6'h00);
        10'h2F9: sin_wave = `S6_TO_U8(6'h00);
        10'h2FA: sin_wave = `S6_TO_U8(6'h00);
        10'h2FB: sin_wave = `S6_TO_U8(6'h00);
        10'h2FC: sin_wave = `S6_TO_U8(6'h00);
        10'h2FD: sin_wave = `S6_TO_U8(6'h00);
        10'h2FE: sin_wave = `S6_TO_U8(6'h00);
        10'h2FF: sin_wave = `S6_TO_U8(6'h00);
        10'h300: sin_wave = `S6_TO_U8(6'h00);
        10'h301: sin_wave = `S6_TO_U8(6'h00);
        10'h302: sin_wave = `S6_TO_U8(6'h00);
        10'h303: sin_wave = `S6_TO_U8(6'h00);
        10'h304: sin_wave = `S6_TO_U8(6'h00);
        10'h305: sin_wave = `S6_TO_U8(6'h00);
        10'h306: sin_wave = `S6_TO_U8(6'h00);
        10'h307: sin_wave = `S6_TO_U8(6'h00);
        10'h308: sin_wave = `S6_TO_U8(6'h00);
        10'h309: sin_wave = `S6_TO_U8(6'h00);
        10'h30A: sin_wave = `S6_TO_U8(6'h00);
        10'h30B: sin_wave = `S6_TO_U8(6'h00);
        10'h30C: sin_wave = `S6_TO_U8(6'h00);
        10'h30D: sin_wave = `S6_TO_U8(6'h00);
        10'h30E: sin_wave = `S6_TO_U8(6'h00);
        10'h30F: sin_wave = `S6_TO_U8(6'h00);
        10'h310: sin_wave = `S6_TO_U8(6'h00);
        10'h311: sin_wave = `S6_TO_U8(6'h00);
        10'h312: sin_wave = `S6_TO_U8(6'h00);
        10'h313: sin_wave = `S6_TO_U8(6'h00);
        10'h314: sin_wave = `S6_TO_U8(6'h00);
        10'h315: sin_wave = `S6_TO_U8(6'h00);
        10'h316: sin_wave = `S6_TO_U8(6'h00);
        10'h317: sin_wave = `S6_TO_U8(6'h00);
        10'h318: sin_wave = `S6_TO_U8(6'h00);
        10'h319: sin_wave = `S6_TO_U8(6'h00);
        10'h31A: sin_wave = `S6_TO_U8(6'h00);
        10'h31B: sin_wave = `S6_TO_U8(6'h00);
        10'h31C: sin_wave = `S6_TO_U8(6'h00);
        10'h31D: sin_wave = `S6_TO_U8(6'h00);
        10'h31E: sin_wave = `S6_TO_U8(6'h00);
        10'h31F: sin_wave = `S6_TO_U8(6'h00);
        10'h320: sin_wave = `S6_TO_U8(6'h00);
        10'h321: sin_wave = `S6_TO_U8(6'h00);
        10'h322: sin_wave = `S6_TO_U8(6'h00);
        10'h323: sin_wave = `S6_TO_U8(6'h00);
        10'h324: sin_wave = `S6_TO_U8(6'h00);
        10'h325: sin_wave = `S6_TO_U8(6'h00);
        10'h326: sin_wave = `S6_TO_U8(6'h00);
        10'h327: sin_wave = `S6_TO_U8(6'h00);
        10'h328: sin_wave = `S6_TO_U8(6'h00);
        10'h329: sin_wave = `S6_TO_U8(6'h00);
        10'h32A: sin_wave = `S6_TO_U8(6'h01);
        10'h32B: sin_wave = `S6_TO_U8(6'h01);
        10'h32C: sin_wave = `S6_TO_U8(6'h01);
        10'h32D: sin_wave = `S6_TO_U8(6'h01);
        10'h32E: sin_wave = `S6_TO_U8(6'h01);
        10'h32F: sin_wave = `S6_TO_U8(6'h01);
        10'h330: sin_wave = `S6_TO_U8(6'h01);
        10'h331: sin_wave = `S6_TO_U8(6'h01);
        10'h332: sin_wave = `S6_TO_U8(6'h01);
        10'h333: sin_wave = `S6_TO_U8(6'h01);
        10'h334: sin_wave = `S6_TO_U8(6'h01);
        10'h335: sin_wave = `S6_TO_U8(6'h01);
        10'h336: sin_wave = `S6_TO_U8(6'h01);
        10'h337: sin_wave = `S6_TO_U8(6'h01);
        10'h338: sin_wave = `S6_TO_U8(6'h01);
        10'h339: sin_wave = `S6_TO_U8(6'h01);
        10'h33A: sin_wave = `S6_TO_U8(6'h01);
        10'h33B: sin_wave = `S6_TO_U8(6'h02);
        10'h33C: sin_wave = `S6_TO_U8(6'h02);
        10'h33D: sin_wave = `S6_TO_U8(6'h02);
        10'h33E: sin_wave = `S6_TO_U8(6'h02);
        10'h33F: sin_wave = `S6_TO_U8(6'h02);
        10'h340: sin_wave = `S6_TO_U8(6'h02);
        10'h341: sin_wave = `S6_TO_U8(6'h02);
        10'h342: sin_wave = `S6_TO_U8(6'h02);
        10'h343: sin_wave = `S6_TO_U8(6'h02);
        10'h344: sin_wave = `S6_TO_U8(6'h02);
        10'h345: sin_wave = `S6_TO_U8(6'h02);
        10'h346: sin_wave = `S6_TO_U8(6'h02);
        10'h347: sin_wave = `S6_TO_U8(6'h02);
        10'h348: sin_wave = `S6_TO_U8(6'h03);
        10'h349: sin_wave = `S6_TO_U8(6'h03);
        10'h34A: sin_wave = `S6_TO_U8(6'h03);
        10'h34B: sin_wave = `S6_TO_U8(6'h03);
        10'h34C: sin_wave = `S6_TO_U8(6'h03);
        10'h34D: sin_wave = `S6_TO_U8(6'h03);
        10'h34E: sin_wave = `S6_TO_U8(6'h03);
        10'h34F: sin_wave = `S6_TO_U8(6'h03);
        10'h350: sin_wave = `S6_TO_U8(6'h03);
        10'h351: sin_wave = `S6_TO_U8(6'h03);
        10'h352: sin_wave = `S6_TO_U8(6'h03);
        10'h353: sin_wave = `S6_TO_U8(6'h03);
        10'h354: sin_wave = `S6_TO_U8(6'h04);
        10'h355: sin_wave = `S6_TO_U8(6'h04);
        10'h356: sin_wave = `S6_TO_U8(6'h04);
        10'h357: sin_wave = `S6_TO_U8(6'h04);
        10'h358: sin_wave = `S6_TO_U8(6'h04);
        10'h359: sin_wave = `S6_TO_U8(6'h04);
        10'h35A: sin_wave = `S6_TO_U8(6'h04);
        10'h35B: sin_wave = `S6_TO_U8(6'h04);
        10'h35C: sin_wave = `S6_TO_U8(6'h04);
        10'h35D: sin_wave = `S6_TO_U8(6'h04);
        10'h35E: sin_wave = `S6_TO_U8(6'h05);
        10'h35F: sin_wave = `S6_TO_U8(6'h05);
        10'h360: sin_wave = `S6_TO_U8(6'h05);
        10'h361: sin_wave = `S6_TO_U8(6'h05);
        10'h362: sin_wave = `S6_TO_U8(6'h05);
        10'h363: sin_wave = `S6_TO_U8(6'h05);
        10'h364: sin_wave = `S6_TO_U8(6'h05);
        10'h365: sin_wave = `S6_TO_U8(6'h05);
        10'h366: sin_wave = `S6_TO_U8(6'h05);
        10'h367: sin_wave = `S6_TO_U8(6'h06);
        10'h368: sin_wave = `S6_TO_U8(6'h06);
        10'h369: sin_wave = `S6_TO_U8(6'h06);
        10'h36A: sin_wave = `S6_TO_U8(6'h06);
        10'h36B: sin_wave = `S6_TO_U8(6'h06);
        10'h36C: sin_wave = `S6_TO_U8(6'h06);
        10'h36D: sin_wave = `S6_TO_U8(6'h06);
        10'h36E: sin_wave = `S6_TO_U8(6'h06);
        10'h36F: sin_wave = `S6_TO_U8(6'h07);
        10'h370: sin_wave = `S6_TO_U8(6'h07);
        10'h371: sin_wave = `S6_TO_U8(6'h07);
        10'h372: sin_wave = `S6_TO_U8(6'h07);
        10'h373: sin_wave = `S6_TO_U8(6'h07);
        10'h374: sin_wave = `S6_TO_U8(6'h07);
        10'h375: sin_wave = `S6_TO_U8(6'h07);
        10'h376: sin_wave = `S6_TO_U8(6'h07);
        10'h377: sin_wave = `S6_TO_U8(6'h08);
        10'h378: sin_wave = `S6_TO_U8(6'h08);
        10'h379: sin_wave = `S6_TO_U8(6'h08);
        10'h37A: sin_wave = `S6_TO_U8(6'h08);
        10'h37B: sin_wave = `S6_TO_U8(6'h08);
        10'h37C: sin_wave = `S6_TO_U8(6'h08);
        10'h37D: sin_wave = `S6_TO_U8(6'h08);
        10'h37E: sin_wave = `S6_TO_U8(6'h08);
        10'h37F: sin_wave = `S6_TO_U8(6'h09);
        10'h380: sin_wave = `S6_TO_U8(6'h09);
        10'h381: sin_wave = `S6_TO_U8(6'h09);
        10'h382: sin_wave = `S6_TO_U8(6'h09);
        10'h383: sin_wave = `S6_TO_U8(6'h09);
        10'h384: sin_wave = `S6_TO_U8(6'h09);
        10'h385: sin_wave = `S6_TO_U8(6'h09);
        10'h386: sin_wave = `S6_TO_U8(6'h0A);
        10'h387: sin_wave = `S6_TO_U8(6'h0A);
        10'h388: sin_wave = `S6_TO_U8(6'h0A);
        10'h389: sin_wave = `S6_TO_U8(6'h0A);
        10'h38A: sin_wave = `S6_TO_U8(6'h0A);
        10'h38B: sin_wave = `S6_TO_U8(6'h0A);
        10'h38C: sin_wave = `S6_TO_U8(6'h0A);
        10'h38D: sin_wave = `S6_TO_U8(6'h0B);
        10'h38E: sin_wave = `S6_TO_U8(6'h0B);
        10'h38F: sin_wave = `S6_TO_U8(6'h0B);
        10'h390: sin_wave = `S6_TO_U8(6'h0B);
        10'h391: sin_wave = `S6_TO_U8(6'h0B);
        10'h392: sin_wave = `S6_TO_U8(6'h0B);
        10'h393: sin_wave = `S6_TO_U8(6'h0B);
        10'h394: sin_wave = `S6_TO_U8(6'h0C);
        10'h395: sin_wave = `S6_TO_U8(6'h0C);
        10'h396: sin_wave = `S6_TO_U8(6'h0C);
        10'h397: sin_wave = `S6_TO_U8(6'h0C);
        10'h398: sin_wave = `S6_TO_U8(6'h0C);
        10'h399: sin_wave = `S6_TO_U8(6'h0C);
        10'h39A: sin_wave = `S6_TO_U8(6'h0D);
        10'h39B: sin_wave = `S6_TO_U8(6'h0D);
        10'h39C: sin_wave = `S6_TO_U8(6'h0D);
        10'h39D: sin_wave = `S6_TO_U8(6'h0D);
        10'h39E: sin_wave = `S6_TO_U8(6'h0D);
        10'h39F: sin_wave = `S6_TO_U8(6'h0D);
        10'h3A0: sin_wave = `S6_TO_U8(6'h0D);
        10'h3A1: sin_wave = `S6_TO_U8(6'h0E);
        10'h3A2: sin_wave = `S6_TO_U8(6'h0E);
        10'h3A3: sin_wave = `S6_TO_U8(6'h0E);
        10'h3A4: sin_wave = `S6_TO_U8(6'h0E);
        10'h3A5: sin_wave = `S6_TO_U8(6'h0E);
        10'h3A6: sin_wave = `S6_TO_U8(6'h0E);
        10'h3A7: sin_wave = `S6_TO_U8(6'h0F);
        10'h3A8: sin_wave = `S6_TO_U8(6'h0F);
        10'h3A9: sin_wave = `S6_TO_U8(6'h0F);
        10'h3AA: sin_wave = `S6_TO_U8(6'h0F);
        10'h3AB: sin_wave = `S6_TO_U8(6'h0F);
        10'h3AC: sin_wave = `S6_TO_U8(6'h0F);
        10'h3AD: sin_wave = `S6_TO_U8(6'h10);
        10'h3AE: sin_wave = `S6_TO_U8(6'h10);
        10'h3AF: sin_wave = `S6_TO_U8(6'h10);
        10'h3B0: sin_wave = `S6_TO_U8(6'h10);
        10'h3B1: sin_wave = `S6_TO_U8(6'h10);
        10'h3B2: sin_wave = `S6_TO_U8(6'h10);
        10'h3B3: sin_wave = `S6_TO_U8(6'h11);
        10'h3B4: sin_wave = `S6_TO_U8(6'h11);
        10'h3B5: sin_wave = `S6_TO_U8(6'h11);
        10'h3B6: sin_wave = `S6_TO_U8(6'h11);
        10'h3B7: sin_wave = `S6_TO_U8(6'h11);
        10'h3B8: sin_wave = `S6_TO_U8(6'h12);
        10'h3B9: sin_wave = `S6_TO_U8(6'h12);
        10'h3BA: sin_wave = `S6_TO_U8(6'h12);
        10'h3BB: sin_wave = `S6_TO_U8(6'h12);
        10'h3BC: sin_wave = `S6_TO_U8(6'h12);
        10'h3BD: sin_wave = `S6_TO_U8(6'h12);
        10'h3BE: sin_wave = `S6_TO_U8(6'h13);
        10'h3BF: sin_wave = `S6_TO_U8(6'h13);
        10'h3C0: sin_wave = `S6_TO_U8(6'h13);
        10'h3C1: sin_wave = `S6_TO_U8(6'h13);
        10'h3C2: sin_wave = `S6_TO_U8(6'h13);
        10'h3C3: sin_wave = `S6_TO_U8(6'h13);
        10'h3C4: sin_wave = `S6_TO_U8(6'h14);
        10'h3C5: sin_wave = `S6_TO_U8(6'h14);
        10'h3C6: sin_wave = `S6_TO_U8(6'h14);
        10'h3C7: sin_wave = `S6_TO_U8(6'h14);
        10'h3C8: sin_wave = `S6_TO_U8(6'h14);
        10'h3C9: sin_wave = `S6_TO_U8(6'h15);
        10'h3CA: sin_wave = `S6_TO_U8(6'h15);
        10'h3CB: sin_wave = `S6_TO_U8(6'h15);
        10'h3CC: sin_wave = `S6_TO_U8(6'h15);
        10'h3CD: sin_wave = `S6_TO_U8(6'h15);
        10'h3CE: sin_wave = `S6_TO_U8(6'h15);
        10'h3CF: sin_wave = `S6_TO_U8(6'h16);
        10'h3D0: sin_wave = `S6_TO_U8(6'h16);
        10'h3D1: sin_wave = `S6_TO_U8(6'h16);
        10'h3D2: sin_wave = `S6_TO_U8(6'h16);
        10'h3D3: sin_wave = `S6_TO_U8(6'h16);
        10'h3D4: sin_wave = `S6_TO_U8(6'h17);
        10'h3D5: sin_wave = `S6_TO_U8(6'h17);
        10'h3D6: sin_wave = `S6_TO_U8(6'h17);
        10'h3D7: sin_wave = `S6_TO_U8(6'h17);
        10'h3D8: sin_wave = `S6_TO_U8(6'h17);
        10'h3D9: sin_wave = `S6_TO_U8(6'h18);
        10'h3DA: sin_wave = `S6_TO_U8(6'h18);
        10'h3DB: sin_wave = `S6_TO_U8(6'h18);
        10'h3DC: sin_wave = `S6_TO_U8(6'h18);
        10'h3DD: sin_wave = `S6_TO_U8(6'h18);
        10'h3DE: sin_wave = `S6_TO_U8(6'h18);
        10'h3DF: sin_wave = `S6_TO_U8(6'h19);
        10'h3E0: sin_wave = `S6_TO_U8(6'h19);
        10'h3E1: sin_wave = `S6_TO_U8(6'h19);
        10'h3E2: sin_wave = `S6_TO_U8(6'h19);
        10'h3E3: sin_wave = `S6_TO_U8(6'h19);
        10'h3E4: sin_wave = `S6_TO_U8(6'h1A);
        10'h3E5: sin_wave = `S6_TO_U8(6'h1A);
        10'h3E6: sin_wave = `S6_TO_U8(6'h1A);
        10'h3E7: sin_wave = `S6_TO_U8(6'h1A);
        10'h3E8: sin_wave = `S6_TO_U8(6'h1A);
        10'h3E9: sin_wave = `S6_TO_U8(6'h1B);
        10'h3EA: sin_wave = `S6_TO_U8(6'h1B);
        10'h3EB: sin_wave = `S6_TO_U8(6'h1B);
        10'h3EC: sin_wave = `S6_TO_U8(6'h1B);
        10'h3ED: sin_wave = `S6_TO_U8(6'h1B);
        10'h3EE: sin_wave = `S6_TO_U8(6'h1C);
        10'h3EF: sin_wave = `S6_TO_U8(6'h1C);
        10'h3F0: sin_wave = `S6_TO_U8(6'h1C);
        10'h3F1: sin_wave = `S6_TO_U8(6'h1C);
        10'h3F2: sin_wave = `S6_TO_U8(6'h1C);
        10'h3F3: sin_wave = `S6_TO_U8(6'h1C);
        10'h3F4: sin_wave = `S6_TO_U8(6'h1D);
        10'h3F5: sin_wave = `S6_TO_U8(6'h1D);
        10'h3F6: sin_wave = `S6_TO_U8(6'h1D);
        10'h3F7: sin_wave = `S6_TO_U8(6'h1D);
        10'h3F8: sin_wave = `S6_TO_U8(6'h1D);
        10'h3F9: sin_wave = `S6_TO_U8(6'h1E);
        10'h3FA: sin_wave = `S6_TO_U8(6'h1E);
        10'h3FB: sin_wave = `S6_TO_U8(6'h1E);
        10'h3FC: sin_wave = `S6_TO_U8(6'h1E);
        10'h3FD: sin_wave = `S6_TO_U8(6'h1E);
        10'h3FE: sin_wave = `S6_TO_U8(6'h1F);
        10'h3FF: sin_wave = `S6_TO_U8(6'h1F);

        default: sin_wave = `S6_TO_U8(6'h00);
    endcase
end

endmodule